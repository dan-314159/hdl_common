module spi_slave(
    );

endmodule
